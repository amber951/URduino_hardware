

 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /xilinx_ram_65536_tb/status
      waveform add -signals /xilinx_ram_65536_tb/xilinx_ram_65536_synth_inst/bmg_port/RSTA
      waveform add -signals /xilinx_ram_65536_tb/xilinx_ram_65536_synth_inst/bmg_port/CLKA
      waveform add -signals /xilinx_ram_65536_tb/xilinx_ram_65536_synth_inst/bmg_port/ADDRA
      waveform add -signals /xilinx_ram_65536_tb/xilinx_ram_65536_synth_inst/bmg_port/DINA
      waveform add -signals /xilinx_ram_65536_tb/xilinx_ram_65536_synth_inst/bmg_port/WEA
      waveform add -signals /xilinx_ram_65536_tb/xilinx_ram_65536_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
